library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity fancy_counter is
    port (
        
    );
end fancy_counter;

architecture Behavioral of fancy_counter is

begin


end Behavioral;
